class transaction;
  rand bit [2:0] a;
  rand bit [2:0] b;
  bit [2:0] y;
endclass