interface and_intf();
  logic [2:0] a;
  logic [2:0] b;
  logic [2:0] y;
endinterface
